library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; -- we need a conversion to unsigned
use WORK.constants.all;

--THE SUM GENERATOR IS ONE OF THE SUB-BLOCKS OF THE PENTIUM 4 ADDER.
--IT IS MADE UP OF SEVERAL CARRY SELECT BLOCKS (#CS-BLOCK = NBIT/NBIT_PER_BLOCK)

--EACH CARRY SELECT BLOCK OPERATES ON A SMALL GROUP OF BITS OF THE TWO OPERANDS
--A AND B (NBIT_PER_BLOCK), COMPUTING THE SUM AMONG THEM.
--EACH BLOCK CALCULATES THE SUM ASSUMING BOTH Cin=0 AND Cin=1 AND THEN IT USES
--THE EFFECTIVE CARRY GENERATED BY THE CARRY GENERATOR TO SELECT THE CORRECT RESULT.


entity SUM_GEN_N is
  generic ( NBIT_PER_BLOCK: integer := numBit;
            NBLOCKS:	integer := 8);
  port (
         A:	in	std_logic_vector(NBIT_PER_BLOCK*NBLOCKS-1 downto 0);
         B:	in	std_logic_vector(NBIT_PER_BLOCK*NBLOCKS-1 downto 0);
         Ci:	in	std_logic_vector(NBLOCKS-1 downto 0);
         S:	out	std_logic_vector(NBIT_PER_BLOCK*NBLOCKS-1 downto 0));
end SUM_GEN_N;


architecture STRUCTURAL of SUM_GEN_N is
  
  component CARRY_SEL_N    
    generic(NBIT: integer := numBit);
    port (A:       in   std_logic_vector(NBIT-1 downto 0);
          B:       in   std_logic_vector(NBIT-1 downto 0);
          Ci:      in   std_logic;
          S:       out  std_logic_vector(NBIT-1 downto 0));
  end component;

  begin

    FOR1: for i in 1 to NBLOCKS generate
      for all: CARRY_SEL_N use configuration WORK.CFG_CARRY_SEL_N;
      begin
        
        UCSi: CARRY_SEL_N
          generic map(NBIT_PER_BLOCK)
          port map (A(i*NBIT_PER_BLOCK-1 downto (i-1)*NBIT_PER_BLOCK), B(i*NBIT_PER_BLOCK-1 downto (i-1)*NBIT_PER_BLOCK), Ci(i-1), S(i*NBIT_PER_BLOCK-1 downto (i-1)*NBIT_PER_BLOCK));
        
    end generate;
    
end STRUCTURAL;

configuration CFG_SUM_GEN_N of SUM_GEN_N is
  for STRUCTURAL
  end for;
end CFG_SUM_GEN_N;
