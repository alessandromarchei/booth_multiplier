library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; -- we need a conversion to unsigned
use WORK.constants.all;

--THE CARRY SELECT ADDER IS MADE UP OF TWO IDENTICAL ADDERS (RCA), EACH GENERATING
--A SET OF SUM BITS AND A CARRY OUT. ACTUALLY, IN THE P4 CARRY SELECT ADDER WE'LL NEGLECT THE CARRY OUT.
--THE TWO ADDERS GENERATE IN PARALLEL THE RESULTS, AS SOON AS INPUTS (A and B)ARRIVES: THE FIRST ONE ASSUMES
--THAT THE INCOMING CARRY IN IS '0', GENERATING THE SUM S0, WHILE THE SECOND ADDER ASSUMES
--THAT THE CARRY IN IS '1', GENERATING THE SUM S1. THE ACTUAL SUM (S) IS SELECTED BY A
--MUX 2 TO 1, WHICH RECIEVES THE EFFECTIVE CARRY IN (Ci) AS SELECTOR SIGNAL.

entity CARRY_SEL_N is
  generic(NBIT: integer := numBit);
  port (A:       in std_logic_vector(NBIT-1 downto 0);
        B:       in std_logic_vector(NBIT-1 downto 0);
        Ci:      in  std_logic;
        S:       out  std_logic_vector(NBIT-1 downto 0));
end CARRY_SEL_N;

architecture STRUCTURAL of CARRY_SEL_N is

  --Declaration of components
  
  component RCAN
        generic ( NBIT : integer := numBit;
                  DRCAS : Time := 0 ns;
	          DRCAC : Time := 0 ns);
	Port (	A:	In	std_logic_vector(NBIT-1 downto 0);
		B:	In	std_logic_vector(NBIT-1 downto 0);
		Ci:	In	std_logic;
		S:	Out	std_logic_vector(NBIT-1 downto 0);
		Co:	Out	std_logic);
  end component;

  component MUX21_GENERIC is
        Generic (NBIT: integer:= numBit;
		 DELAY_MUX: Time:= tp_mux);
	Port (	A:	In	std_logic_vector(NBIT-1 downto 0);
                B:	In	std_logic_vector(NBIT-1 downto 0);
		SEL:	In	std_logic;
		Y:	Out	std_logic_vector(NBIT-1 downto 0));
  end component;

  signal S1, S0: std_logic_vector(NBIT-1 downto 0);
  signal Cout0, Cout1: std_logic; --signals containing the useless carry out generated by the two
                                  --adders
                                              
  begin

     RCA1: RCAN 
	   generic map (NBIT, DRCAS => 0.2 ns, DRCAC => 0.2 ns)
           port map (A, B, '1', S1, Cout1);
     
     RCA0: RCAN 
	   generic map (NBIT, DRCAS => 0.2 ns, DRCAC => 0.2 ns)
           port map (A, B, '0', S0, Cout0);

     MUX21: MUX21_GENERIC
	   generic map (NBIT, DELAY_MUX => 0.5 ns )
	   port map (S0, S1, Ci, S);

    
end STRUCTURAL;

configuration CFG_CARRY_SEL_N of CARRY_SEL_N is
  
  for STRUCTURAL
    
    for RCA1: RCAN
      use configuration WORK.CFG_RCAN_STRUCTURAL;
    end for;
    
    for RCA0: RCAN
      use configuration WORK.CFG_RCAN_STRUCTURAL;
    end for;
    
    for MUX21: MUX21_GENERIC
      use configuration WORK.CFG_MUX21_GEN_STRUCTURAL;
    end for;
    
  end for;
  
end CFG_CARRY_SEL_N;
