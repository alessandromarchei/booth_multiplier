library IEEE;
use IEEE.std_logic_1164.all; --  libreria IEEE con definizione tipi standard logic
use WORK.constants.all; -- libreria WORK user-defined


--THIS MODULE HAS BEEN DESIGNED IN ORDER TO IMPLEMENT THE BOOTH'S ALGORITHM.

--BY EXTRACTING A TRIPLET OF BITS FROM THE MULTIPLIER IT IS ABLE TO GENERATE A
--TRIPLET OF BITS TO SELECT PROPERLY THE INPUT OF A 5 TO 1 MUX WHICH
--CORRESPONDS TO THE PARTIAL SUM OF THE ALGORITHM.

--THE OUTPUT OF OUR ENCODER WILL BE THEN CONNECTED TO THE SELECTOR OF THE
--MODULE CALLED "MUX51_GENERIC" INSIDE THE HIGHER LEVEL DESIGN CALLED "BOOTHMUL".

entity ENCODER is
	Port (	INPUT:	In	std_logic_vector(2 downto 0) ;
		OUTPUT: Out	std_logic_vector(2 downto 0));
end ENCODER;


architecture BEHAVIORAL of ENCODER is

-- FROM THE TRUTH TABLE WE FOUND THE RELATIONSHIPS AMONG THE TRIPLET AT THE
-- INPUT AND FOR EACH BIT OF THE OUTPUT TRIPLET

--THIS WAY WE TRIED TO OPTIMIZE AGAIN THE IMPLEMENTATION OF THE CIRCUIT,
--INSTEAD OF USING A BEHAVIORAL APPROACH THAT COULD RESULT IN A MORE GENERIC BEHAVIOR
begin
  --LSB of the output
out0 : OUTPUT(0) <= (not(INPUT(2)) and INPUT(0)) or (not(INPUT(2)) and INPUT(1));

out1 : OUTPUT(1) <= (not(INPUT(2)) and INPUT(1) and INPUT(0)) or (INPUT(2) and (NOT(INPUT(1))) and INPUT(0)) or (INPUT(2) and INPUT(1) and (NOT(INPUT(0))));

  --MSB OF THE OUTPUT
out2 : OUTPUT(2) <= INPUT(2) and (NOT(INPUT(1))) and (NOT(INPUT(0)));             

end BEHAVIORAL;



